
//`timescale 1ps/1ps

module tb_top;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
endmodule

