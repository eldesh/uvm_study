`include "sample_seq_item.sv"
`include "sample_master_seq_lib.sv"
`include "sample_slave_seq_lib.sv"
`include "sample_scrbd_item.sv"

`include "sample_master_driver.sv"
`include "sample_master_monitor.sv"
`include "sample_master_sequencer.sv"
`include "sample_master_agent.sv"

`include "sample_slave_driver.sv"
`include "sample_slave_sequencer.sv"
`include "sample_slave_agent.sv"

`include "sample_env.sv"
